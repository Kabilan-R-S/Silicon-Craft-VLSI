module hello();
  initial
    $display("HELLO WORLD");
endmodule
